// layer_encoding.vh
//
// Copyright (C) 2020 Dan Rodrigues <danrr.gh.oss@gmail.com>
//
// SPDX-License-Identifier: Apache-2.0

`ifndef layer_encoding_vh
`define layer_encoding_vh

`define LAYER_SPRITES 4
`define LAYER_SCROLL3 3
`define LAYER_SCROLL2 2
`define LAYER_SCROLL1 1
`define LAYER_SCROLL0 0

`define LAYER_SPRITES_OHE (1 << 4)
`define LAYER_SCROLL3_OHE (1 << 3)
`define LAYER_SCROLL2_OHE (1 << 2)
`define LAYER_SCROLL1_OHE (1 << 1)
`define LAYER_SCROLL0_OHE (1 << 0)

`endif
