VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vdp_lite_user_proj
  CLASS BLOCK ;
  FOREIGN vdp_lite_user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 1400.000 BY 1100.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 1096.000 274.530 1100.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 261.160 1400.000 261.760 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.610 1096.000 1132.890 1100.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 1096.000 344.450 1100.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.050 1096.000 909.330 1100.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.530 0.000 1110.810 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.010 1096.000 714.290 1100.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 54.440 1400.000 55.040 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1111.450 1096.000 1111.730 1100.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.970 0.000 1209.250 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 786.120 1400.000 786.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 1096.000 163.210 1100.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 706.650 1096.000 706.930 1100.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.770 1096.000 763.050 1100.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.050 1096.000 679.330 1100.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 817.400 1400.000 818.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1362.610 1096.000 1362.890 1100.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 497.800 1400.000 498.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1054.040 1400.000 1054.640 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.890 1096.000 888.170 1100.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 1096.000 316.850 1100.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.210 1096.000 470.490 1100.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 486.920 1400.000 487.520 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 930.280 1400.000 930.880 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 342.760 1400.000 343.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 1096.000 484.290 1100.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.930 0.000 1313.210 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 322.360 1400.000 322.960 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 532.770 1096.000 533.050 1100.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 909.880 1400.000 910.480 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1096.000 1062.970 1100.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1074.440 1400.000 1075.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1285.330 1096.000 1285.610 1100.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.250 0.000 1125.530 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 1096.000 860.570 1100.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 1096.000 309.490 1100.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.250 1096.000 205.530 1100.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.010 1096.000 254.290 1100.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 538.600 1400.000 539.200 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1341.450 1096.000 1341.730 1100.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 574.170 1096.000 574.450 1100.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1396.650 1096.000 1396.930 1100.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1174.010 1096.000 1174.290 1100.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.250 1096.000 504.530 1100.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.050 1096.000 449.330 1100.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 457.000 1400.000 457.600 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 961.560 1400.000 962.160 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 1096.000 79.490 1100.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 936.650 1096.000 936.930 1100.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 569.880 1400.000 570.480 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1044.520 4.000 1045.120 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 1096.000 511.890 1100.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1013.240 1400.000 1013.840 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.970 1096.000 749.250 1100.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1382.850 0.000 1383.130 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 965.170 1096.000 965.450 1100.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.210 1096.000 700.490 1100.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.090 1096.000 414.370 1100.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 44.920 1400.000 45.520 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 992.840 1400.000 993.440 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 985.410 1096.000 985.690 1100.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 209.480 1400.000 210.080 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.610 1096.000 1201.890 1100.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.530 1096.000 351.810 1100.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1361.690 0.000 1361.970 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.530 1096.000 581.810 1100.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1265.090 1096.000 1265.370 1100.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.570 1096.000 1006.850 1100.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 126.520 1400.000 127.120 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.090 1096.000 1334.370 1100.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 595.330 1096.000 595.610 1100.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.650 1096.000 1097.930 1100.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 1096.000 211.970 1100.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 1096.000 30.730 1100.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 291.080 1400.000 291.680 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 776.600 1400.000 777.200 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 1096.000 246.930 1100.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1085.320 1400.000 1085.920 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 671.690 1096.000 671.970 1100.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.450 1096.000 490.730 1100.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 1096.000 1195.450 1100.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 34.040 1400.000 34.640 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 972.440 1400.000 973.040 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 425.720 1400.000 426.320 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 631.080 1400.000 631.680 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.130 1096.000 609.410 1100.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 23.160 1400.000 23.760 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.370 1096.000 560.650 1100.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 961.560 4.000 962.160 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1002.360 1400.000 1002.960 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 301.960 1400.000 302.560 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 754.840 1400.000 755.440 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.530 1096.000 1041.810 1100.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 1096.000 24.290 1100.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 1096.000 142.050 1100.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 848.680 1400.000 849.280 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 693.640 1400.000 694.240 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 1096.000 44.530 1100.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.010 1096.000 944.290 1100.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.970 1096.000 128.250 1100.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.810 1096.000 958.090 1100.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 1096.000 198.170 1100.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 1096.000 1055.610 1100.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 724.920 1400.000 725.520 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 405.320 1400.000 405.920 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.290 1096.000 1090.570 1100.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1347.890 1096.000 1348.170 1100.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 941.160 1400.000 941.760 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 981.960 1400.000 982.560 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.770 0.000 1062.050 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1117.890 1096.000 1118.170 1100.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.730 0.000 1258.010 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 4.000 869.680 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.930 1096.000 1083.210 1100.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 270.680 1400.000 271.280 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.130 1096.000 149.410 1100.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1033.640 1400.000 1034.240 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.450 1096.000 950.730 1100.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 1096.000 289.250 1100.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.250 1096.000 435.530 1100.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 189.080 1400.000 189.680 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1306.490 0.000 1306.770 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.730 0.000 1097.010 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 529.080 1400.000 529.680 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 950.680 1400.000 951.280 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.410 1096.000 755.690 1100.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 1096.000 86.850 1100.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.810 1096.000 498.090 1100.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.450 1096.000 651.730 1100.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1230.130 1096.000 1230.410 1100.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 427.890 1096.000 428.170 1100.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 13.640 1400.000 14.240 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 1096.000 16.930 1100.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 559.000 1400.000 559.600 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1117.890 0.000 1118.170 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 374.040 1400.000 374.640 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 1096.000 93.290 1100.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 1096.000 65.690 1100.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 1096.000 38.090 1100.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1313.850 1096.000 1314.130 1100.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.490 1096.000 225.770 1100.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1257.730 1096.000 1258.010 1100.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1022.760 1400.000 1023.360 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 198.600 1400.000 199.200 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 363.160 1400.000 363.760 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 665.250 1096.000 665.530 1100.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 371.770 1096.000 372.050 1100.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.730 1096.000 1028.010 1100.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1396.650 0.000 1396.930 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.530 0.000 1041.810 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 895.250 1096.000 895.530 1100.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1000.130 1096.000 1000.410 1100.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.050 0.000 1139.330 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 525.410 1096.000 525.690 1100.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 745.320 1400.000 745.920 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.170 1096.000 804.450 1100.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 869.080 1400.000 869.680 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.210 1096.000 539.490 1100.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 146.920 1400.000 147.520 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 920.760 1400.000 921.360 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 508.680 1400.000 509.280 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 250.280 1400.000 250.880 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 239.400 1400.000 240.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1104.090 1096.000 1104.370 1100.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1222.770 0.000 1223.050 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 65.320 1400.000 65.920 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 673.240 1400.000 673.840 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 337.730 1096.000 338.010 1100.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 1096.000 190.810 1100.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 1096.000 1146.690 1100.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.130 1096.000 1069.410 1100.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 518.200 1400.000 518.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.930 1096.000 623.210 1100.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 811.530 1096.000 811.810 1100.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1382.850 1096.000 1383.130 1100.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 386.490 1096.000 386.770 1100.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 1096.000 114.450 1100.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 837.800 1400.000 838.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1208.970 1096.000 1209.250 1100.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.970 1096.000 979.250 1100.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 167.320 1400.000 167.920 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 765.720 1400.000 766.320 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 922.850 1096.000 923.130 1100.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 394.440 1400.000 395.040 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.250 1096.000 1125.530 1100.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.930 1096.000 784.210 1100.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 414.840 1400.000 415.440 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 602.690 1096.000 602.970 1100.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1355.250 1096.000 1355.530 1100.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 85.720 1400.000 86.320 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1166.650 1096.000 1166.930 1100.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 446.120 1400.000 446.720 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 1096.000 3.130 1100.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 1096.000 135.610 1100.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.730 1096.000 177.010 1100.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 353.640 1400.000 354.240 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.290 1096.000 630.570 1100.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 333.240 1400.000 333.840 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 1096.000 379.410 1100.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1320.290 1096.000 1320.570 1100.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1278.890 1096.000 1279.170 1100.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 1096.000 233.130 1100.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 734.440 1400.000 735.040 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 797.730 1096.000 798.010 1100.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 477.400 1400.000 478.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 281.560 1400.000 282.160 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 797.000 1400.000 797.600 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 735.170 1096.000 735.450 1100.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 590.280 1400.000 590.880 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.610 1096.000 741.890 1100.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.890 1096.000 1049.170 1100.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.330 0.000 825.610 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 1096.000 121.810 1100.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 1096.000 588.250 1100.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 1096.000 853.210 1100.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 95.240 1400.000 95.840 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.970 1096.000 519.250 1100.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1096.000 1014.210 1100.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1044.520 1400.000 1045.120 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1347.890 0.000 1348.170 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1181.370 1096.000 1181.650 1100.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 106.120 1400.000 106.720 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 157.800 1400.000 158.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 714.040 1400.000 714.640 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 901.690 1096.000 901.970 1100.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 435.240 1400.000 435.840 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.450 1096.000 881.730 1100.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1375.490 0.000 1375.770 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 662.360 1400.000 662.960 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.410 0.000 1215.690 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 1096.000 463.130 1100.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 1096.000 365.610 1100.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.290 1096.000 239.570 1100.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.720 4.000 1004.320 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 682.760 1400.000 683.360 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 878.600 1400.000 879.200 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.370 1096.000 1250.650 1100.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 704.520 1400.000 705.120 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 1096.000 170.570 1100.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.690 0.000 1292.970 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.410 1096.000 1215.690 1100.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 621.560 1400.000 622.160 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 178.200 1400.000 178.800 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 832.690 1096.000 832.970 1100.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 916.410 1096.000 916.690 1100.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.730 1096.000 637.010 1100.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.810 1096.000 1188.090 1100.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 549.480 1400.000 550.080 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.450 1096.000 421.730 1100.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.050 1096.000 1369.330 1100.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.290 1096.000 400.570 1100.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.490 1096.000 1076.770 1100.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 1096.000 51.890 1100.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 826.920 1400.000 827.520 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.690 1096.000 441.970 1100.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 1096.000 58.330 1100.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 1096.000 776.850 1100.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 229.880 1400.000 230.480 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.530 1096.000 1271.810 1100.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 900.360 1400.000 900.960 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 1096.000 73.050 1100.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1034.170 1096.000 1034.450 1100.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1236.570 1096.000 1236.850 1100.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 1096.000 107.090 1100.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 117.000 1400.000 117.600 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 476.650 1096.000 476.930 1100.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.330 1096.000 825.610 1100.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 610.680 1400.000 611.280 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.930 1096.000 393.210 1100.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 1096.000 100.650 1100.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.450 1096.000 260.730 1100.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.050 0.000 1369.330 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.210 1096.000 930.490 1100.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 137.400 1400.000 138.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 806.520 1400.000 807.120 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.410 1096.000 1376.690 1100.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.960 4.000 982.560 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.490 1096.000 685.770 1100.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.090 0.000 1334.370 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1096.000 1153.130 1100.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 992.770 1096.000 993.050 1100.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 1096.000 184.370 1100.000 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 692.850 1096.000 693.130 1100.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 889.480 1400.000 890.080 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.010 1096.000 323.290 1100.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.050 1096.000 219.330 1100.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.490 1096.000 846.770 1100.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 1096.000 281.890 1100.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.690 1096.000 1292.970 1100.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 1096.000 1020.650 1100.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 74.840 1400.000 75.440 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.370 1096.000 790.650 1100.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1327.650 1096.000 1327.930 1100.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 652.840 1400.000 653.440 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.210 1096.000 769.490 1100.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.930 1096.000 554.210 1100.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 641.960 1400.000 642.560 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.970 1096.000 818.250 1100.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 219.000 1400.000 219.600 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.810 1096.000 728.090 1100.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.970 1096.000 358.250 1100.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1306.490 1096.000 1306.770 1100.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 1096.000 1299.410 1100.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1064.920 1400.000 1065.520 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 1096.000 1160.490 1100.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 1096.000 330.650 1100.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 1096.000 9.570 1100.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 1096.000 867.930 1100.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 580.760 1400.000 581.360 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 601.160 1400.000 601.760 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 295.410 1096.000 295.690 1100.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1355.250 0.000 1355.530 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.810 0.000 958.090 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 466.520 1400.000 467.120 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.090 1096.000 874.370 1100.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.890 1096.000 658.170 1100.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.770 1096.000 1223.050 1100.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 1096.000 720.730 1100.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.770 1096.000 303.050 1100.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1390.210 1096.000 1390.490 1100.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1243.930 1096.000 1244.210 1100.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 1096.000 455.770 1100.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.490 1096.000 616.770 1100.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.570 1096.000 546.850 1100.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 858.200 1400.000 858.800 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.090 1096.000 644.370 1100.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.810 1096.000 268.090 1100.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.730 1096.000 568.010 1100.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.050 1096.000 1139.330 1100.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 971.610 1096.000 971.890 1100.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.730 1096.000 407.010 1100.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 1096.000 156.770 1100.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 384.920 1400.000 385.520 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 839.130 1096.000 839.410 1100.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 312.840 1400.000 313.440 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1394.260 1088.085 ;
      LAYER met1 ;
        RECT 2.830 4.460 1396.950 1095.780 ;
      LAYER met2 ;
        RECT 3.410 1095.720 9.010 1096.000 ;
        RECT 9.850 1095.720 16.370 1096.000 ;
        RECT 17.210 1095.720 23.730 1096.000 ;
        RECT 24.570 1095.720 30.170 1096.000 ;
        RECT 31.010 1095.720 37.530 1096.000 ;
        RECT 38.370 1095.720 43.970 1096.000 ;
        RECT 44.810 1095.720 51.330 1096.000 ;
        RECT 52.170 1095.720 57.770 1096.000 ;
        RECT 58.610 1095.720 65.130 1096.000 ;
        RECT 65.970 1095.720 72.490 1096.000 ;
        RECT 73.330 1095.720 78.930 1096.000 ;
        RECT 79.770 1095.720 86.290 1096.000 ;
        RECT 87.130 1095.720 92.730 1096.000 ;
        RECT 93.570 1095.720 100.090 1096.000 ;
        RECT 100.930 1095.720 106.530 1096.000 ;
        RECT 107.370 1095.720 113.890 1096.000 ;
        RECT 114.730 1095.720 121.250 1096.000 ;
        RECT 122.090 1095.720 127.690 1096.000 ;
        RECT 128.530 1095.720 135.050 1096.000 ;
        RECT 135.890 1095.720 141.490 1096.000 ;
        RECT 142.330 1095.720 148.850 1096.000 ;
        RECT 149.690 1095.720 156.210 1096.000 ;
        RECT 157.050 1095.720 162.650 1096.000 ;
        RECT 163.490 1095.720 170.010 1096.000 ;
        RECT 170.850 1095.720 176.450 1096.000 ;
        RECT 177.290 1095.720 183.810 1096.000 ;
        RECT 184.650 1095.720 190.250 1096.000 ;
        RECT 191.090 1095.720 197.610 1096.000 ;
        RECT 198.450 1095.720 204.970 1096.000 ;
        RECT 205.810 1095.720 211.410 1096.000 ;
        RECT 212.250 1095.720 218.770 1096.000 ;
        RECT 219.610 1095.720 225.210 1096.000 ;
        RECT 226.050 1095.720 232.570 1096.000 ;
        RECT 233.410 1095.720 239.010 1096.000 ;
        RECT 239.850 1095.720 246.370 1096.000 ;
        RECT 247.210 1095.720 253.730 1096.000 ;
        RECT 254.570 1095.720 260.170 1096.000 ;
        RECT 261.010 1095.720 267.530 1096.000 ;
        RECT 268.370 1095.720 273.970 1096.000 ;
        RECT 274.810 1095.720 281.330 1096.000 ;
        RECT 282.170 1095.720 288.690 1096.000 ;
        RECT 289.530 1095.720 295.130 1096.000 ;
        RECT 295.970 1095.720 302.490 1096.000 ;
        RECT 303.330 1095.720 308.930 1096.000 ;
        RECT 309.770 1095.720 316.290 1096.000 ;
        RECT 317.130 1095.720 322.730 1096.000 ;
        RECT 323.570 1095.720 330.090 1096.000 ;
        RECT 330.930 1095.720 337.450 1096.000 ;
        RECT 338.290 1095.720 343.890 1096.000 ;
        RECT 344.730 1095.720 351.250 1096.000 ;
        RECT 352.090 1095.720 357.690 1096.000 ;
        RECT 358.530 1095.720 365.050 1096.000 ;
        RECT 365.890 1095.720 371.490 1096.000 ;
        RECT 372.330 1095.720 378.850 1096.000 ;
        RECT 379.690 1095.720 386.210 1096.000 ;
        RECT 387.050 1095.720 392.650 1096.000 ;
        RECT 393.490 1095.720 400.010 1096.000 ;
        RECT 400.850 1095.720 406.450 1096.000 ;
        RECT 407.290 1095.720 413.810 1096.000 ;
        RECT 414.650 1095.720 421.170 1096.000 ;
        RECT 422.010 1095.720 427.610 1096.000 ;
        RECT 428.450 1095.720 434.970 1096.000 ;
        RECT 435.810 1095.720 441.410 1096.000 ;
        RECT 442.250 1095.720 448.770 1096.000 ;
        RECT 449.610 1095.720 455.210 1096.000 ;
        RECT 456.050 1095.720 462.570 1096.000 ;
        RECT 463.410 1095.720 469.930 1096.000 ;
        RECT 470.770 1095.720 476.370 1096.000 ;
        RECT 477.210 1095.720 483.730 1096.000 ;
        RECT 484.570 1095.720 490.170 1096.000 ;
        RECT 491.010 1095.720 497.530 1096.000 ;
        RECT 498.370 1095.720 503.970 1096.000 ;
        RECT 504.810 1095.720 511.330 1096.000 ;
        RECT 512.170 1095.720 518.690 1096.000 ;
        RECT 519.530 1095.720 525.130 1096.000 ;
        RECT 525.970 1095.720 532.490 1096.000 ;
        RECT 533.330 1095.720 538.930 1096.000 ;
        RECT 539.770 1095.720 546.290 1096.000 ;
        RECT 547.130 1095.720 553.650 1096.000 ;
        RECT 554.490 1095.720 560.090 1096.000 ;
        RECT 560.930 1095.720 567.450 1096.000 ;
        RECT 568.290 1095.720 573.890 1096.000 ;
        RECT 574.730 1095.720 581.250 1096.000 ;
        RECT 582.090 1095.720 587.690 1096.000 ;
        RECT 588.530 1095.720 595.050 1096.000 ;
        RECT 595.890 1095.720 602.410 1096.000 ;
        RECT 603.250 1095.720 608.850 1096.000 ;
        RECT 609.690 1095.720 616.210 1096.000 ;
        RECT 617.050 1095.720 622.650 1096.000 ;
        RECT 623.490 1095.720 630.010 1096.000 ;
        RECT 630.850 1095.720 636.450 1096.000 ;
        RECT 637.290 1095.720 643.810 1096.000 ;
        RECT 644.650 1095.720 651.170 1096.000 ;
        RECT 652.010 1095.720 657.610 1096.000 ;
        RECT 658.450 1095.720 664.970 1096.000 ;
        RECT 665.810 1095.720 671.410 1096.000 ;
        RECT 672.250 1095.720 678.770 1096.000 ;
        RECT 679.610 1095.720 685.210 1096.000 ;
        RECT 686.050 1095.720 692.570 1096.000 ;
        RECT 693.410 1095.720 699.930 1096.000 ;
        RECT 700.770 1095.720 706.370 1096.000 ;
        RECT 707.210 1095.720 713.730 1096.000 ;
        RECT 714.570 1095.720 720.170 1096.000 ;
        RECT 721.010 1095.720 727.530 1096.000 ;
        RECT 728.370 1095.720 734.890 1096.000 ;
        RECT 735.730 1095.720 741.330 1096.000 ;
        RECT 742.170 1095.720 748.690 1096.000 ;
        RECT 749.530 1095.720 755.130 1096.000 ;
        RECT 755.970 1095.720 762.490 1096.000 ;
        RECT 763.330 1095.720 768.930 1096.000 ;
        RECT 769.770 1095.720 776.290 1096.000 ;
        RECT 777.130 1095.720 783.650 1096.000 ;
        RECT 784.490 1095.720 790.090 1096.000 ;
        RECT 790.930 1095.720 797.450 1096.000 ;
        RECT 798.290 1095.720 803.890 1096.000 ;
        RECT 804.730 1095.720 811.250 1096.000 ;
        RECT 812.090 1095.720 817.690 1096.000 ;
        RECT 818.530 1095.720 825.050 1096.000 ;
        RECT 825.890 1095.720 832.410 1096.000 ;
        RECT 833.250 1095.720 838.850 1096.000 ;
        RECT 839.690 1095.720 846.210 1096.000 ;
        RECT 847.050 1095.720 852.650 1096.000 ;
        RECT 853.490 1095.720 860.010 1096.000 ;
        RECT 860.850 1095.720 867.370 1096.000 ;
        RECT 868.210 1095.720 873.810 1096.000 ;
        RECT 874.650 1095.720 881.170 1096.000 ;
        RECT 882.010 1095.720 887.610 1096.000 ;
        RECT 888.450 1095.720 894.970 1096.000 ;
        RECT 895.810 1095.720 901.410 1096.000 ;
        RECT 902.250 1095.720 908.770 1096.000 ;
        RECT 909.610 1095.720 916.130 1096.000 ;
        RECT 916.970 1095.720 922.570 1096.000 ;
        RECT 923.410 1095.720 929.930 1096.000 ;
        RECT 930.770 1095.720 936.370 1096.000 ;
        RECT 937.210 1095.720 943.730 1096.000 ;
        RECT 944.570 1095.720 950.170 1096.000 ;
        RECT 951.010 1095.720 957.530 1096.000 ;
        RECT 958.370 1095.720 964.890 1096.000 ;
        RECT 965.730 1095.720 971.330 1096.000 ;
        RECT 972.170 1095.720 978.690 1096.000 ;
        RECT 979.530 1095.720 985.130 1096.000 ;
        RECT 985.970 1095.720 992.490 1096.000 ;
        RECT 993.330 1095.720 999.850 1096.000 ;
        RECT 1000.690 1095.720 1006.290 1096.000 ;
        RECT 1007.130 1095.720 1013.650 1096.000 ;
        RECT 1014.490 1095.720 1020.090 1096.000 ;
        RECT 1020.930 1095.720 1027.450 1096.000 ;
        RECT 1028.290 1095.720 1033.890 1096.000 ;
        RECT 1034.730 1095.720 1041.250 1096.000 ;
        RECT 1042.090 1095.720 1048.610 1096.000 ;
        RECT 1049.450 1095.720 1055.050 1096.000 ;
        RECT 1055.890 1095.720 1062.410 1096.000 ;
        RECT 1063.250 1095.720 1068.850 1096.000 ;
        RECT 1069.690 1095.720 1076.210 1096.000 ;
        RECT 1077.050 1095.720 1082.650 1096.000 ;
        RECT 1083.490 1095.720 1090.010 1096.000 ;
        RECT 1090.850 1095.720 1097.370 1096.000 ;
        RECT 1098.210 1095.720 1103.810 1096.000 ;
        RECT 1104.650 1095.720 1111.170 1096.000 ;
        RECT 1112.010 1095.720 1117.610 1096.000 ;
        RECT 1118.450 1095.720 1124.970 1096.000 ;
        RECT 1125.810 1095.720 1132.330 1096.000 ;
        RECT 1133.170 1095.720 1138.770 1096.000 ;
        RECT 1139.610 1095.720 1146.130 1096.000 ;
        RECT 1146.970 1095.720 1152.570 1096.000 ;
        RECT 1153.410 1095.720 1159.930 1096.000 ;
        RECT 1160.770 1095.720 1166.370 1096.000 ;
        RECT 1167.210 1095.720 1173.730 1096.000 ;
        RECT 1174.570 1095.720 1181.090 1096.000 ;
        RECT 1181.930 1095.720 1187.530 1096.000 ;
        RECT 1188.370 1095.720 1194.890 1096.000 ;
        RECT 1195.730 1095.720 1201.330 1096.000 ;
        RECT 1202.170 1095.720 1208.690 1096.000 ;
        RECT 1209.530 1095.720 1215.130 1096.000 ;
        RECT 1215.970 1095.720 1222.490 1096.000 ;
        RECT 1223.330 1095.720 1229.850 1096.000 ;
        RECT 1230.690 1095.720 1236.290 1096.000 ;
        RECT 1237.130 1095.720 1243.650 1096.000 ;
        RECT 1244.490 1095.720 1250.090 1096.000 ;
        RECT 1250.930 1095.720 1257.450 1096.000 ;
        RECT 1258.290 1095.720 1264.810 1096.000 ;
        RECT 1265.650 1095.720 1271.250 1096.000 ;
        RECT 1272.090 1095.720 1278.610 1096.000 ;
        RECT 1279.450 1095.720 1285.050 1096.000 ;
        RECT 1285.890 1095.720 1292.410 1096.000 ;
        RECT 1293.250 1095.720 1298.850 1096.000 ;
        RECT 1299.690 1095.720 1306.210 1096.000 ;
        RECT 1307.050 1095.720 1313.570 1096.000 ;
        RECT 1314.410 1095.720 1320.010 1096.000 ;
        RECT 1320.850 1095.720 1327.370 1096.000 ;
        RECT 1328.210 1095.720 1333.810 1096.000 ;
        RECT 1334.650 1095.720 1341.170 1096.000 ;
        RECT 1342.010 1095.720 1347.610 1096.000 ;
        RECT 1348.450 1095.720 1354.970 1096.000 ;
        RECT 1355.810 1095.720 1362.330 1096.000 ;
        RECT 1363.170 1095.720 1368.770 1096.000 ;
        RECT 1369.610 1095.720 1376.130 1096.000 ;
        RECT 1376.970 1095.720 1382.570 1096.000 ;
        RECT 1383.410 1095.720 1389.930 1096.000 ;
        RECT 1390.770 1095.720 1396.370 1096.000 ;
        RECT 2.860 4.280 1396.920 1095.720 ;
        RECT 3.410 4.000 9.010 4.280 ;
        RECT 9.850 4.000 16.370 4.280 ;
        RECT 17.210 4.000 22.810 4.280 ;
        RECT 23.650 4.000 30.170 4.280 ;
        RECT 31.010 4.000 36.610 4.280 ;
        RECT 37.450 4.000 43.970 4.280 ;
        RECT 44.810 4.000 51.330 4.280 ;
        RECT 52.170 4.000 57.770 4.280 ;
        RECT 58.610 4.000 65.130 4.280 ;
        RECT 65.970 4.000 71.570 4.280 ;
        RECT 72.410 4.000 78.930 4.280 ;
        RECT 79.770 4.000 85.370 4.280 ;
        RECT 86.210 4.000 92.730 4.280 ;
        RECT 93.570 4.000 100.090 4.280 ;
        RECT 100.930 4.000 106.530 4.280 ;
        RECT 107.370 4.000 113.890 4.280 ;
        RECT 114.730 4.000 120.330 4.280 ;
        RECT 121.170 4.000 127.690 4.280 ;
        RECT 128.530 4.000 134.130 4.280 ;
        RECT 134.970 4.000 141.490 4.280 ;
        RECT 142.330 4.000 148.850 4.280 ;
        RECT 149.690 4.000 155.290 4.280 ;
        RECT 156.130 4.000 162.650 4.280 ;
        RECT 163.490 4.000 169.090 4.280 ;
        RECT 169.930 4.000 176.450 4.280 ;
        RECT 177.290 4.000 183.810 4.280 ;
        RECT 184.650 4.000 190.250 4.280 ;
        RECT 191.090 4.000 197.610 4.280 ;
        RECT 198.450 4.000 204.050 4.280 ;
        RECT 204.890 4.000 211.410 4.280 ;
        RECT 212.250 4.000 217.850 4.280 ;
        RECT 218.690 4.000 225.210 4.280 ;
        RECT 226.050 4.000 232.570 4.280 ;
        RECT 233.410 4.000 239.010 4.280 ;
        RECT 239.850 4.000 246.370 4.280 ;
        RECT 247.210 4.000 252.810 4.280 ;
        RECT 253.650 4.000 260.170 4.280 ;
        RECT 261.010 4.000 266.610 4.280 ;
        RECT 267.450 4.000 273.970 4.280 ;
        RECT 274.810 4.000 281.330 4.280 ;
        RECT 282.170 4.000 287.770 4.280 ;
        RECT 288.610 4.000 295.130 4.280 ;
        RECT 295.970 4.000 301.570 4.280 ;
        RECT 302.410 4.000 308.930 4.280 ;
        RECT 309.770 4.000 316.290 4.280 ;
        RECT 317.130 4.000 322.730 4.280 ;
        RECT 323.570 4.000 330.090 4.280 ;
        RECT 330.930 4.000 336.530 4.280 ;
        RECT 337.370 4.000 343.890 4.280 ;
        RECT 344.730 4.000 350.330 4.280 ;
        RECT 351.170 4.000 357.690 4.280 ;
        RECT 358.530 4.000 365.050 4.280 ;
        RECT 365.890 4.000 371.490 4.280 ;
        RECT 372.330 4.000 378.850 4.280 ;
        RECT 379.690 4.000 385.290 4.280 ;
        RECT 386.130 4.000 392.650 4.280 ;
        RECT 393.490 4.000 399.090 4.280 ;
        RECT 399.930 4.000 406.450 4.280 ;
        RECT 407.290 4.000 413.810 4.280 ;
        RECT 414.650 4.000 420.250 4.280 ;
        RECT 421.090 4.000 427.610 4.280 ;
        RECT 428.450 4.000 434.050 4.280 ;
        RECT 434.890 4.000 441.410 4.280 ;
        RECT 442.250 4.000 448.770 4.280 ;
        RECT 449.610 4.000 455.210 4.280 ;
        RECT 456.050 4.000 462.570 4.280 ;
        RECT 463.410 4.000 469.010 4.280 ;
        RECT 469.850 4.000 476.370 4.280 ;
        RECT 477.210 4.000 482.810 4.280 ;
        RECT 483.650 4.000 490.170 4.280 ;
        RECT 491.010 4.000 497.530 4.280 ;
        RECT 498.370 4.000 503.970 4.280 ;
        RECT 504.810 4.000 511.330 4.280 ;
        RECT 512.170 4.000 517.770 4.280 ;
        RECT 518.610 4.000 525.130 4.280 ;
        RECT 525.970 4.000 531.570 4.280 ;
        RECT 532.410 4.000 538.930 4.280 ;
        RECT 539.770 4.000 546.290 4.280 ;
        RECT 547.130 4.000 552.730 4.280 ;
        RECT 553.570 4.000 560.090 4.280 ;
        RECT 560.930 4.000 566.530 4.280 ;
        RECT 567.370 4.000 573.890 4.280 ;
        RECT 574.730 4.000 581.250 4.280 ;
        RECT 582.090 4.000 587.690 4.280 ;
        RECT 588.530 4.000 595.050 4.280 ;
        RECT 595.890 4.000 601.490 4.280 ;
        RECT 602.330 4.000 608.850 4.280 ;
        RECT 609.690 4.000 615.290 4.280 ;
        RECT 616.130 4.000 622.650 4.280 ;
        RECT 623.490 4.000 630.010 4.280 ;
        RECT 630.850 4.000 636.450 4.280 ;
        RECT 637.290 4.000 643.810 4.280 ;
        RECT 644.650 4.000 650.250 4.280 ;
        RECT 651.090 4.000 657.610 4.280 ;
        RECT 658.450 4.000 664.050 4.280 ;
        RECT 664.890 4.000 671.410 4.280 ;
        RECT 672.250 4.000 678.770 4.280 ;
        RECT 679.610 4.000 685.210 4.280 ;
        RECT 686.050 4.000 692.570 4.280 ;
        RECT 693.410 4.000 699.010 4.280 ;
        RECT 699.850 4.000 706.370 4.280 ;
        RECT 707.210 4.000 713.730 4.280 ;
        RECT 714.570 4.000 720.170 4.280 ;
        RECT 721.010 4.000 727.530 4.280 ;
        RECT 728.370 4.000 733.970 4.280 ;
        RECT 734.810 4.000 741.330 4.280 ;
        RECT 742.170 4.000 747.770 4.280 ;
        RECT 748.610 4.000 755.130 4.280 ;
        RECT 755.970 4.000 762.490 4.280 ;
        RECT 763.330 4.000 768.930 4.280 ;
        RECT 769.770 4.000 776.290 4.280 ;
        RECT 777.130 4.000 782.730 4.280 ;
        RECT 783.570 4.000 790.090 4.280 ;
        RECT 790.930 4.000 796.530 4.280 ;
        RECT 797.370 4.000 803.890 4.280 ;
        RECT 804.730 4.000 811.250 4.280 ;
        RECT 812.090 4.000 817.690 4.280 ;
        RECT 818.530 4.000 825.050 4.280 ;
        RECT 825.890 4.000 831.490 4.280 ;
        RECT 832.330 4.000 838.850 4.280 ;
        RECT 839.690 4.000 845.290 4.280 ;
        RECT 846.130 4.000 852.650 4.280 ;
        RECT 853.490 4.000 860.010 4.280 ;
        RECT 860.850 4.000 866.450 4.280 ;
        RECT 867.290 4.000 873.810 4.280 ;
        RECT 874.650 4.000 880.250 4.280 ;
        RECT 881.090 4.000 887.610 4.280 ;
        RECT 888.450 4.000 894.970 4.280 ;
        RECT 895.810 4.000 901.410 4.280 ;
        RECT 902.250 4.000 908.770 4.280 ;
        RECT 909.610 4.000 915.210 4.280 ;
        RECT 916.050 4.000 922.570 4.280 ;
        RECT 923.410 4.000 929.010 4.280 ;
        RECT 929.850 4.000 936.370 4.280 ;
        RECT 937.210 4.000 943.730 4.280 ;
        RECT 944.570 4.000 950.170 4.280 ;
        RECT 951.010 4.000 957.530 4.280 ;
        RECT 958.370 4.000 963.970 4.280 ;
        RECT 964.810 4.000 971.330 4.280 ;
        RECT 972.170 4.000 977.770 4.280 ;
        RECT 978.610 4.000 985.130 4.280 ;
        RECT 985.970 4.000 992.490 4.280 ;
        RECT 993.330 4.000 998.930 4.280 ;
        RECT 999.770 4.000 1006.290 4.280 ;
        RECT 1007.130 4.000 1012.730 4.280 ;
        RECT 1013.570 4.000 1020.090 4.280 ;
        RECT 1020.930 4.000 1027.450 4.280 ;
        RECT 1028.290 4.000 1033.890 4.280 ;
        RECT 1034.730 4.000 1041.250 4.280 ;
        RECT 1042.090 4.000 1047.690 4.280 ;
        RECT 1048.530 4.000 1055.050 4.280 ;
        RECT 1055.890 4.000 1061.490 4.280 ;
        RECT 1062.330 4.000 1068.850 4.280 ;
        RECT 1069.690 4.000 1076.210 4.280 ;
        RECT 1077.050 4.000 1082.650 4.280 ;
        RECT 1083.490 4.000 1090.010 4.280 ;
        RECT 1090.850 4.000 1096.450 4.280 ;
        RECT 1097.290 4.000 1103.810 4.280 ;
        RECT 1104.650 4.000 1110.250 4.280 ;
        RECT 1111.090 4.000 1117.610 4.280 ;
        RECT 1118.450 4.000 1124.970 4.280 ;
        RECT 1125.810 4.000 1131.410 4.280 ;
        RECT 1132.250 4.000 1138.770 4.280 ;
        RECT 1139.610 4.000 1145.210 4.280 ;
        RECT 1146.050 4.000 1152.570 4.280 ;
        RECT 1153.410 4.000 1159.930 4.280 ;
        RECT 1160.770 4.000 1166.370 4.280 ;
        RECT 1167.210 4.000 1173.730 4.280 ;
        RECT 1174.570 4.000 1180.170 4.280 ;
        RECT 1181.010 4.000 1187.530 4.280 ;
        RECT 1188.370 4.000 1193.970 4.280 ;
        RECT 1194.810 4.000 1201.330 4.280 ;
        RECT 1202.170 4.000 1208.690 4.280 ;
        RECT 1209.530 4.000 1215.130 4.280 ;
        RECT 1215.970 4.000 1222.490 4.280 ;
        RECT 1223.330 4.000 1228.930 4.280 ;
        RECT 1229.770 4.000 1236.290 4.280 ;
        RECT 1237.130 4.000 1242.730 4.280 ;
        RECT 1243.570 4.000 1250.090 4.280 ;
        RECT 1250.930 4.000 1257.450 4.280 ;
        RECT 1258.290 4.000 1263.890 4.280 ;
        RECT 1264.730 4.000 1271.250 4.280 ;
        RECT 1272.090 4.000 1277.690 4.280 ;
        RECT 1278.530 4.000 1285.050 4.280 ;
        RECT 1285.890 4.000 1292.410 4.280 ;
        RECT 1293.250 4.000 1298.850 4.280 ;
        RECT 1299.690 4.000 1306.210 4.280 ;
        RECT 1307.050 4.000 1312.650 4.280 ;
        RECT 1313.490 4.000 1320.010 4.280 ;
        RECT 1320.850 4.000 1326.450 4.280 ;
        RECT 1327.290 4.000 1333.810 4.280 ;
        RECT 1334.650 4.000 1341.170 4.280 ;
        RECT 1342.010 4.000 1347.610 4.280 ;
        RECT 1348.450 4.000 1354.970 4.280 ;
        RECT 1355.810 4.000 1361.410 4.280 ;
        RECT 1362.250 4.000 1368.770 4.280 ;
        RECT 1369.610 4.000 1375.210 4.280 ;
        RECT 1376.050 4.000 1382.570 4.280 ;
        RECT 1383.410 4.000 1389.930 4.280 ;
        RECT 1390.770 4.000 1396.370 4.280 ;
      LAYER met3 ;
        RECT 4.000 1086.320 1396.000 1088.165 ;
        RECT 4.400 1084.920 1395.600 1086.320 ;
        RECT 4.000 1076.800 1396.000 1084.920 ;
        RECT 4.400 1075.440 1396.000 1076.800 ;
        RECT 4.400 1075.400 1395.600 1075.440 ;
        RECT 4.000 1074.040 1395.600 1075.400 ;
        RECT 4.000 1065.920 1396.000 1074.040 ;
        RECT 4.400 1064.520 1395.600 1065.920 ;
        RECT 4.000 1055.040 1396.000 1064.520 ;
        RECT 4.400 1053.640 1395.600 1055.040 ;
        RECT 4.000 1045.520 1396.000 1053.640 ;
        RECT 4.400 1044.120 1395.600 1045.520 ;
        RECT 4.000 1034.640 1396.000 1044.120 ;
        RECT 4.400 1033.240 1395.600 1034.640 ;
        RECT 4.000 1025.120 1396.000 1033.240 ;
        RECT 4.400 1023.760 1396.000 1025.120 ;
        RECT 4.400 1023.720 1395.600 1023.760 ;
        RECT 4.000 1022.360 1395.600 1023.720 ;
        RECT 4.000 1014.240 1396.000 1022.360 ;
        RECT 4.400 1012.840 1395.600 1014.240 ;
        RECT 4.000 1004.720 1396.000 1012.840 ;
        RECT 4.400 1003.360 1396.000 1004.720 ;
        RECT 4.400 1003.320 1395.600 1003.360 ;
        RECT 4.000 1001.960 1395.600 1003.320 ;
        RECT 4.000 993.840 1396.000 1001.960 ;
        RECT 4.400 992.440 1395.600 993.840 ;
        RECT 4.000 982.960 1396.000 992.440 ;
        RECT 4.400 981.560 1395.600 982.960 ;
        RECT 4.000 973.440 1396.000 981.560 ;
        RECT 4.400 972.040 1395.600 973.440 ;
        RECT 4.000 962.560 1396.000 972.040 ;
        RECT 4.400 961.160 1395.600 962.560 ;
        RECT 4.000 953.040 1396.000 961.160 ;
        RECT 4.400 951.680 1396.000 953.040 ;
        RECT 4.400 951.640 1395.600 951.680 ;
        RECT 4.000 950.280 1395.600 951.640 ;
        RECT 4.000 942.160 1396.000 950.280 ;
        RECT 4.400 940.760 1395.600 942.160 ;
        RECT 4.000 932.640 1396.000 940.760 ;
        RECT 4.400 931.280 1396.000 932.640 ;
        RECT 4.400 931.240 1395.600 931.280 ;
        RECT 4.000 929.880 1395.600 931.240 ;
        RECT 4.000 921.760 1396.000 929.880 ;
        RECT 4.400 920.360 1395.600 921.760 ;
        RECT 4.000 910.880 1396.000 920.360 ;
        RECT 4.400 909.480 1395.600 910.880 ;
        RECT 4.000 901.360 1396.000 909.480 ;
        RECT 4.400 899.960 1395.600 901.360 ;
        RECT 4.000 890.480 1396.000 899.960 ;
        RECT 4.400 889.080 1395.600 890.480 ;
        RECT 4.000 880.960 1396.000 889.080 ;
        RECT 4.400 879.600 1396.000 880.960 ;
        RECT 4.400 879.560 1395.600 879.600 ;
        RECT 4.000 878.200 1395.600 879.560 ;
        RECT 4.000 870.080 1396.000 878.200 ;
        RECT 4.400 868.680 1395.600 870.080 ;
        RECT 4.000 860.560 1396.000 868.680 ;
        RECT 4.400 859.200 1396.000 860.560 ;
        RECT 4.400 859.160 1395.600 859.200 ;
        RECT 4.000 857.800 1395.600 859.160 ;
        RECT 4.000 849.680 1396.000 857.800 ;
        RECT 4.400 848.280 1395.600 849.680 ;
        RECT 4.000 838.800 1396.000 848.280 ;
        RECT 4.400 837.400 1395.600 838.800 ;
        RECT 4.000 829.280 1396.000 837.400 ;
        RECT 4.400 827.920 1396.000 829.280 ;
        RECT 4.400 827.880 1395.600 827.920 ;
        RECT 4.000 826.520 1395.600 827.880 ;
        RECT 4.000 818.400 1396.000 826.520 ;
        RECT 4.400 817.000 1395.600 818.400 ;
        RECT 4.000 808.880 1396.000 817.000 ;
        RECT 4.400 807.520 1396.000 808.880 ;
        RECT 4.400 807.480 1395.600 807.520 ;
        RECT 4.000 806.120 1395.600 807.480 ;
        RECT 4.000 798.000 1396.000 806.120 ;
        RECT 4.400 796.600 1395.600 798.000 ;
        RECT 4.000 787.120 1396.000 796.600 ;
        RECT 4.400 785.720 1395.600 787.120 ;
        RECT 4.000 777.600 1396.000 785.720 ;
        RECT 4.400 776.200 1395.600 777.600 ;
        RECT 4.000 766.720 1396.000 776.200 ;
        RECT 4.400 765.320 1395.600 766.720 ;
        RECT 4.000 757.200 1396.000 765.320 ;
        RECT 4.400 755.840 1396.000 757.200 ;
        RECT 4.400 755.800 1395.600 755.840 ;
        RECT 4.000 754.440 1395.600 755.800 ;
        RECT 4.000 746.320 1396.000 754.440 ;
        RECT 4.400 744.920 1395.600 746.320 ;
        RECT 4.000 736.800 1396.000 744.920 ;
        RECT 4.400 735.440 1396.000 736.800 ;
        RECT 4.400 735.400 1395.600 735.440 ;
        RECT 4.000 734.040 1395.600 735.400 ;
        RECT 4.000 725.920 1396.000 734.040 ;
        RECT 4.400 724.520 1395.600 725.920 ;
        RECT 4.000 715.040 1396.000 724.520 ;
        RECT 4.400 713.640 1395.600 715.040 ;
        RECT 4.000 705.520 1396.000 713.640 ;
        RECT 4.400 704.120 1395.600 705.520 ;
        RECT 4.000 694.640 1396.000 704.120 ;
        RECT 4.400 693.240 1395.600 694.640 ;
        RECT 4.000 685.120 1396.000 693.240 ;
        RECT 4.400 683.760 1396.000 685.120 ;
        RECT 4.400 683.720 1395.600 683.760 ;
        RECT 4.000 682.360 1395.600 683.720 ;
        RECT 4.000 674.240 1396.000 682.360 ;
        RECT 4.400 672.840 1395.600 674.240 ;
        RECT 4.000 664.720 1396.000 672.840 ;
        RECT 4.400 663.360 1396.000 664.720 ;
        RECT 4.400 663.320 1395.600 663.360 ;
        RECT 4.000 661.960 1395.600 663.320 ;
        RECT 4.000 653.840 1396.000 661.960 ;
        RECT 4.400 652.440 1395.600 653.840 ;
        RECT 4.000 642.960 1396.000 652.440 ;
        RECT 4.400 641.560 1395.600 642.960 ;
        RECT 4.000 633.440 1396.000 641.560 ;
        RECT 4.400 632.080 1396.000 633.440 ;
        RECT 4.400 632.040 1395.600 632.080 ;
        RECT 4.000 630.680 1395.600 632.040 ;
        RECT 4.000 622.560 1396.000 630.680 ;
        RECT 4.400 621.160 1395.600 622.560 ;
        RECT 4.000 613.040 1396.000 621.160 ;
        RECT 4.400 611.680 1396.000 613.040 ;
        RECT 4.400 611.640 1395.600 611.680 ;
        RECT 4.000 610.280 1395.600 611.640 ;
        RECT 4.000 602.160 1396.000 610.280 ;
        RECT 4.400 600.760 1395.600 602.160 ;
        RECT 4.000 591.280 1396.000 600.760 ;
        RECT 4.400 589.880 1395.600 591.280 ;
        RECT 4.000 581.760 1396.000 589.880 ;
        RECT 4.400 580.360 1395.600 581.760 ;
        RECT 4.000 570.880 1396.000 580.360 ;
        RECT 4.400 569.480 1395.600 570.880 ;
        RECT 4.000 561.360 1396.000 569.480 ;
        RECT 4.400 560.000 1396.000 561.360 ;
        RECT 4.400 559.960 1395.600 560.000 ;
        RECT 4.000 558.600 1395.600 559.960 ;
        RECT 4.000 550.480 1396.000 558.600 ;
        RECT 4.400 549.080 1395.600 550.480 ;
        RECT 4.000 540.960 1396.000 549.080 ;
        RECT 4.400 539.600 1396.000 540.960 ;
        RECT 4.400 539.560 1395.600 539.600 ;
        RECT 4.000 538.200 1395.600 539.560 ;
        RECT 4.000 530.080 1396.000 538.200 ;
        RECT 4.400 528.680 1395.600 530.080 ;
        RECT 4.000 519.200 1396.000 528.680 ;
        RECT 4.400 517.800 1395.600 519.200 ;
        RECT 4.000 509.680 1396.000 517.800 ;
        RECT 4.400 508.280 1395.600 509.680 ;
        RECT 4.000 498.800 1396.000 508.280 ;
        RECT 4.400 497.400 1395.600 498.800 ;
        RECT 4.000 489.280 1396.000 497.400 ;
        RECT 4.400 487.920 1396.000 489.280 ;
        RECT 4.400 487.880 1395.600 487.920 ;
        RECT 4.000 486.520 1395.600 487.880 ;
        RECT 4.000 478.400 1396.000 486.520 ;
        RECT 4.400 477.000 1395.600 478.400 ;
        RECT 4.000 468.880 1396.000 477.000 ;
        RECT 4.400 467.520 1396.000 468.880 ;
        RECT 4.400 467.480 1395.600 467.520 ;
        RECT 4.000 466.120 1395.600 467.480 ;
        RECT 4.000 458.000 1396.000 466.120 ;
        RECT 4.400 456.600 1395.600 458.000 ;
        RECT 4.000 447.120 1396.000 456.600 ;
        RECT 4.400 445.720 1395.600 447.120 ;
        RECT 4.000 437.600 1396.000 445.720 ;
        RECT 4.400 436.240 1396.000 437.600 ;
        RECT 4.400 436.200 1395.600 436.240 ;
        RECT 4.000 434.840 1395.600 436.200 ;
        RECT 4.000 426.720 1396.000 434.840 ;
        RECT 4.400 425.320 1395.600 426.720 ;
        RECT 4.000 417.200 1396.000 425.320 ;
        RECT 4.400 415.840 1396.000 417.200 ;
        RECT 4.400 415.800 1395.600 415.840 ;
        RECT 4.000 414.440 1395.600 415.800 ;
        RECT 4.000 406.320 1396.000 414.440 ;
        RECT 4.400 404.920 1395.600 406.320 ;
        RECT 4.000 395.440 1396.000 404.920 ;
        RECT 4.400 394.040 1395.600 395.440 ;
        RECT 4.000 385.920 1396.000 394.040 ;
        RECT 4.400 384.520 1395.600 385.920 ;
        RECT 4.000 375.040 1396.000 384.520 ;
        RECT 4.400 373.640 1395.600 375.040 ;
        RECT 4.000 365.520 1396.000 373.640 ;
        RECT 4.400 364.160 1396.000 365.520 ;
        RECT 4.400 364.120 1395.600 364.160 ;
        RECT 4.000 362.760 1395.600 364.120 ;
        RECT 4.000 354.640 1396.000 362.760 ;
        RECT 4.400 353.240 1395.600 354.640 ;
        RECT 4.000 345.120 1396.000 353.240 ;
        RECT 4.400 343.760 1396.000 345.120 ;
        RECT 4.400 343.720 1395.600 343.760 ;
        RECT 4.000 342.360 1395.600 343.720 ;
        RECT 4.000 334.240 1396.000 342.360 ;
        RECT 4.400 332.840 1395.600 334.240 ;
        RECT 4.000 323.360 1396.000 332.840 ;
        RECT 4.400 321.960 1395.600 323.360 ;
        RECT 4.000 313.840 1396.000 321.960 ;
        RECT 4.400 312.440 1395.600 313.840 ;
        RECT 4.000 302.960 1396.000 312.440 ;
        RECT 4.400 301.560 1395.600 302.960 ;
        RECT 4.000 293.440 1396.000 301.560 ;
        RECT 4.400 292.080 1396.000 293.440 ;
        RECT 4.400 292.040 1395.600 292.080 ;
        RECT 4.000 290.680 1395.600 292.040 ;
        RECT 4.000 282.560 1396.000 290.680 ;
        RECT 4.400 281.160 1395.600 282.560 ;
        RECT 4.000 273.040 1396.000 281.160 ;
        RECT 4.400 271.680 1396.000 273.040 ;
        RECT 4.400 271.640 1395.600 271.680 ;
        RECT 4.000 270.280 1395.600 271.640 ;
        RECT 4.000 262.160 1396.000 270.280 ;
        RECT 4.400 260.760 1395.600 262.160 ;
        RECT 4.000 251.280 1396.000 260.760 ;
        RECT 4.400 249.880 1395.600 251.280 ;
        RECT 4.000 241.760 1396.000 249.880 ;
        RECT 4.400 240.400 1396.000 241.760 ;
        RECT 4.400 240.360 1395.600 240.400 ;
        RECT 4.000 239.000 1395.600 240.360 ;
        RECT 4.000 230.880 1396.000 239.000 ;
        RECT 4.400 229.480 1395.600 230.880 ;
        RECT 4.000 221.360 1396.000 229.480 ;
        RECT 4.400 220.000 1396.000 221.360 ;
        RECT 4.400 219.960 1395.600 220.000 ;
        RECT 4.000 218.600 1395.600 219.960 ;
        RECT 4.000 210.480 1396.000 218.600 ;
        RECT 4.400 209.080 1395.600 210.480 ;
        RECT 4.000 199.600 1396.000 209.080 ;
        RECT 4.400 198.200 1395.600 199.600 ;
        RECT 4.000 190.080 1396.000 198.200 ;
        RECT 4.400 188.680 1395.600 190.080 ;
        RECT 4.000 179.200 1396.000 188.680 ;
        RECT 4.400 177.800 1395.600 179.200 ;
        RECT 4.000 169.680 1396.000 177.800 ;
        RECT 4.400 168.320 1396.000 169.680 ;
        RECT 4.400 168.280 1395.600 168.320 ;
        RECT 4.000 166.920 1395.600 168.280 ;
        RECT 4.000 158.800 1396.000 166.920 ;
        RECT 4.400 157.400 1395.600 158.800 ;
        RECT 4.000 149.280 1396.000 157.400 ;
        RECT 4.400 147.920 1396.000 149.280 ;
        RECT 4.400 147.880 1395.600 147.920 ;
        RECT 4.000 146.520 1395.600 147.880 ;
        RECT 4.000 138.400 1396.000 146.520 ;
        RECT 4.400 137.000 1395.600 138.400 ;
        RECT 4.000 127.520 1396.000 137.000 ;
        RECT 4.400 126.120 1395.600 127.520 ;
        RECT 4.000 118.000 1396.000 126.120 ;
        RECT 4.400 116.600 1395.600 118.000 ;
        RECT 4.000 107.120 1396.000 116.600 ;
        RECT 4.400 105.720 1395.600 107.120 ;
        RECT 4.000 97.600 1396.000 105.720 ;
        RECT 4.400 96.240 1396.000 97.600 ;
        RECT 4.400 96.200 1395.600 96.240 ;
        RECT 4.000 94.840 1395.600 96.200 ;
        RECT 4.000 86.720 1396.000 94.840 ;
        RECT 4.400 85.320 1395.600 86.720 ;
        RECT 4.000 77.200 1396.000 85.320 ;
        RECT 4.400 75.840 1396.000 77.200 ;
        RECT 4.400 75.800 1395.600 75.840 ;
        RECT 4.000 74.440 1395.600 75.800 ;
        RECT 4.000 66.320 1396.000 74.440 ;
        RECT 4.400 64.920 1395.600 66.320 ;
        RECT 4.000 55.440 1396.000 64.920 ;
        RECT 4.400 54.040 1395.600 55.440 ;
        RECT 4.000 45.920 1396.000 54.040 ;
        RECT 4.400 44.520 1395.600 45.920 ;
        RECT 4.000 35.040 1396.000 44.520 ;
        RECT 4.400 33.640 1395.600 35.040 ;
        RECT 4.000 25.520 1396.000 33.640 ;
        RECT 4.400 24.160 1396.000 25.520 ;
        RECT 4.400 24.120 1395.600 24.160 ;
        RECT 4.000 22.760 1395.600 24.120 ;
        RECT 4.000 14.640 1396.000 22.760 ;
        RECT 4.400 13.240 1395.600 14.640 ;
        RECT 4.000 10.715 1396.000 13.240 ;
      LAYER met4 ;
        RECT 44.455 10.640 97.440 1088.240 ;
        RECT 99.840 10.640 1328.240 1088.240 ;
  END
END vdp_lite_user_proj
END LIBRARY

